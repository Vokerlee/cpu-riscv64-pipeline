// General data types
`define BYTE_BITS  8
`define HWORD_BITS 16
`define WORD_BITS  32
`define DWORD_BITS 64

// ALU defines
`define ALU_ADD  4'b0000
`define ALU_SUB  4'b0001
`define ALU_AND  4'b0010
`define ALU_OR   4'b0011
`define ALU_XOR  4'b0100
`define ALU_SHL  4'b1000
`define ALU_SHR  4'b1001
`define ALU_SHA  4'b1010
`define ALU_SLT  4'b1011
`define ALU_SLTU 4'b1100
